class Frame;
  
       bit [ 3 :  0] strobe = 4'hF;
       bit [31 :  0] data;
  
endclass