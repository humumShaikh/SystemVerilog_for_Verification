interface intf();

  logic A;
  logic B;
  logic Y;

endinterface