//Basic Interface 
//Just declare all the ports of your DUT

interface intf();

  logic A;
  logic B;
  logic Y;

endinterface
