//Interface (not a class , it is static and not dynamic)
//Just declare all your DUT ports here

interface intf();

  logic A;
  logic B;
  logic Y;

endinterface