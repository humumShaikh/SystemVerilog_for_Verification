interface intf();

  logic A;
  logic B;
  logic [1:0] S;
  logic Y;

endinterface