//Absolutely Basic Interface
//Just define all your DUT ports here , in our case it's a simple 2 input OR Gate
//Declare the ports as type 'logic'

interface intf();

  logic A;    
  logic B;
  logic Y;

endinterface
