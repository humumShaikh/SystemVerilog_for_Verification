//Basic interface 
//Just declare all the ports as 'logic' type that are in your DUT
interface intf();

  logic A;
  logic B;
  logic Y;

endinterface
