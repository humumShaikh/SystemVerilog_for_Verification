//Basic Or-Gate Design File

module orGate
(
  input wire A,
  input wire B,
  output wire Y
);

  assign Y = A | B;

endmodule
